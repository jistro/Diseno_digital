library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
 
entity RljC_Min_U is
    PORT (
        clk    : IN  STD_LOGIC;
        areset : IN  STD_LOGIC;
        aload  : IN  STD_LOGIC;
        data   : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        --cnt_out: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		S0 : OUT  STD_LOGIC;
		S1 : OUT  STD_LOGIC;
		S2 : OUT  STD_LOGIC;
        S3 : OUT  STD_LOGIC;
        UPD: OUT  STD_LOGIC
    );
end RljC_Min_U;
 
architecture Behavioral of RljC_Min_U is
    signal cnt_tmp : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
    signal flag_upd: STD_LOGIC_VECTOR(0 DOWNTO 0) := "0";
begin
    proceso_contador: process (aload, areset, clk, data) begin
        if areset = '1' then
            cnt_tmp <= "0000";
        elsif aload = '1' then
            cnt_tmp <= data;
        elsif rising_edge(clk) then
            if cnt_tmp = "1001" then --cuando detecte reloj a "9"
                cnt_tmp <= "0000";
                flag_upd(0) <= '1';
            else
                cnt_tmp <= cnt_tmp + 1;
                flag_upd(0) <= '0';
            end if;
        end if;
    end process;
	 S0  <= cnt_tmp(0);
	 S1  <= cnt_tmp(1);
	 S2  <= cnt_tmp(2);
     S3  <= cnt_tmp(3);
     UPD <= flag_upd(0);
end Behavioral;
